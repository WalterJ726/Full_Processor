/**
 * NOTE: you should not need to change this file! This file will be swapped out for a grading
 * "skeleton" for testing. We will also remove your imem and dmem file.
 *
 * NOTE: skeleton should be your top-level module!
 *
 * This skeleton file serves as a wrapper around the processor to provide certain control signals
 * and interfaces to memory elements. This structure allows for easier testing, as it is easier to
 * inspect which signals the processor tries to assert when.
 */

module skeleton(clock, reset, imem_clock, dmem_clock, processor_clock, regfile_clock
,address_imem, q_imem, address_dmem, data, wren, q_dmem, ctrl_writeEnable, ctrl_writeReg,
ctrl_readRegA, ctrl_readRegB, data_writeReg, data_readRegA, data_readRegB//, outputWrite
);
    input clock, reset;
    output imem_clock, dmem_clock, processor_clock, regfile_clock;
	 
	 wire clk_div2, clk_div4;
	 frequency_divider frediv_1(clock,reset,clk_div2);
	 frequency_divider frediv_2(clk_div2,reset,clk_div4);
	 assign imem_clock = clock;
	 assign regfile_clock = ~clk_div4;
	 assign processor_clock = ~clk_div4;
	 assign dmem_clock = ~clk_div2;
	 
//	 	wire clk_div2, clk_div4, clk_div8;
//	 frequency_divider frediv_1(clock,reset,clk_div2);
//	 frequency_divider frediv_2(clk_div2,reset,clk_div4);
//	 frequency_divider frediv_3(clk_div4,reset,clk_div8);
//	 assign imem_clock = ~clk_div2;
//	 assign dmem_clock = ~clk_div2;
//	 assign regfile_clock = clk_div4;
//	 assign processor_clock = clk_div8;
    /** IMEM **/
    // Figure out how to generate a Quartus syncram component and commit the generated verilog file.
    // Make sure you configure it correctly!
//    output wire [11:0] address_imem;
//    output wire [31:0] q_imem;
    output [11:0] address_imem;
    output [31:0] q_imem;
    imem my_imem(
        .address    (address_imem),            // address of data
        .clock      (imem_clock),             // you may need to invert the clock
        .q          (q_imem)                   // the raw instruction
    );

    /** DMEM **/
    // Figure out how to generate a Quartus syncram component and commit the generated verilog file.
    // Make sure you configure it correctly!
//    output wire [11:0] address_dmem;
//    output wire [31:0] data;
//    output wire wren;
//    output wire [31:0] q_dmem;
    output [11:0] address_dmem;
    output  [31:0] data;
    output  wren;
    output [31:0] q_dmem;
    dmem my_dmem(
        .address    (address_dmem),       // address of data
        .clock      (dmem_clock),        // may need to invert the clock
        .data	    (data),                // data you want to write
        .wren	    (wren),                // write enable
        .q          (q_dmem)              // data from dmem
    );

    /** REGFILE **/
    // Instantiate your regfile
//    output wire ctrl_writeEnable;
//    output wire [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
//    output wire [31:0] data_writeReg;
//    output wire [31:0] data_readRegA, data_readRegB;
    output ctrl_writeEnable;
    output [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
    output [31:0] data_writeReg;
    output [31:0] data_readRegA, data_readRegB;
	 //output wire [31:0] outputWrite;
    regfile my_regfile(
        regfile_clock,
        ctrl_writeEnable,
        reset,
        ctrl_writeReg,
        ctrl_readRegA,
        ctrl_readRegB,
        data_writeReg,
        data_readRegA,
        data_readRegB
		  //,outputWrite
    );

    /** PROCESSOR **/
    processor my_processor(
        // Control signals
        processor_clock,                // I: The master clock
        reset,                          // I: A reset signal

        // Imem
        address_imem,                   // O: The address of the data to get from imem
        q_imem,                         // I: The data from imem

        // Dmem
        address_dmem,                   // O: The address of the data to get or put from/to dmem
        data,                           // O: The data to write to dmem
        wren,                           // O: Write enable for dmem
        q_dmem,                         // I: The data from dmem

        // Regfile
        ctrl_writeEnable,               // O: Write enable for regfile
        ctrl_writeReg,                  // O: Register to write to in regfile
        ctrl_readRegA,                  // O: Register to read from port A of regfile
        ctrl_readRegB,                  // O: Register to read from port B of regfile
        data_writeReg,                  // O: Data to write to for regfile
        data_readRegA,                  // I: Data from port A of regfile
        data_readRegB                   // I: Data from port B of regfile
    );

endmodule