module extend(ext_immediate,immediate);
	input [16:0] immediate;
	output [31:0] ext_immediate;
	assign ext_immediate[0]=immediate[0];
	assign ext_immediate[1]=immediate[1];
	assign ext_immediate[2]=immediate[2];
	assign ext_immediate[3]=immediate[3];
	assign ext_immediate[4]=immediate[4];
	assign ext_immediate[5]=immediate[5];
	assign ext_immediate[6]=immediate[6];
	assign ext_immediate[7]=immediate[7];
	assign ext_immediate[8]=immediate[8];
	assign ext_immediate[9]=immediate[9];
	assign ext_immediate[10]=immediate[10];
	assign ext_immediate[11]=immediate[11];
	assign ext_immediate[12]=immediate[12];
	assign ext_immediate[13]=immediate[13];
	assign ext_immediate[14]=immediate[14];
	assign ext_immediate[15]=immediate[15];
	assign ext_immediate[16]=immediate[16];
	assign ext_immediate[17]=immediate[16];
	assign ext_immediate[18]=immediate[16];
	assign ext_immediate[19]=immediate[16];
	assign ext_immediate[20]=immediate[16];
	assign ext_immediate[21]=immediate[16];
	assign ext_immediate[22]=immediate[16];
	assign ext_immediate[23]=immediate[16];
	assign ext_immediate[24]=immediate[16];
	assign ext_immediate[25]=immediate[16];
	assign ext_immediate[26]=immediate[16];
	assign ext_immediate[27]=immediate[16];
	assign ext_immediate[28]=immediate[16];
	assign ext_immediate[29]=immediate[16];
	assign ext_immediate[30]=immediate[16];
	assign ext_immediate[31]=immediate[16];
	
	endmodule
	