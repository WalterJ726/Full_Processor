module sra(out,in,shift);
	output [31:0] out;
	input [31:0] in;
	input [4:0] shift;
	
	wire [31:0] out1,out2,out3,out4;
	
	wire most_significant;
	and (most_significant,in[31],1);
	// first layer 1
	assign out1[31] = shift[0] ? most_significant : in[31];
	assign out1[30] = shift[0] ? in[31] : in[30];
	assign out1[29] = shift[0] ? in[30] : in[29];
	assign out1[28] = shift[0] ? in[29] : in[28];
	assign out1[27] = shift[0] ? in[28] : in[27];
	assign out1[26] = shift[0] ? in[27] : in[26];
	assign out1[25] = shift[0] ? in[26] : in[25];
	assign out1[24] = shift[0] ? in[25] : in[24];
	assign out1[23] = shift[0] ? in[24] : in[23];
	assign out1[22] = shift[0] ? in[23] : in[22];
	assign out1[21] = shift[0] ? in[22] : in[21];
	assign out1[20] = shift[0] ? in[21] : in[20];
	assign out1[19] = shift[0] ? in[20] : in[19];
	assign out1[18] = shift[0] ? in[19] : in[18];
	assign out1[17] = shift[0] ? in[18] : in[17];
	assign out1[16] = shift[0] ? in[17] : in[16];
	assign out1[15] = shift[0] ? in[16] : in[15];
	assign out1[14] = shift[0] ? in[15] : in[14];
	assign out1[13] = shift[0] ? in[14] : in[13];
	assign out1[12] = shift[0] ? in[13] : in[12];
	assign out1[11] = shift[0] ? in[12] : in[11];
	assign out1[10] = shift[0] ? in[11] : in[10];
	assign out1[9] = shift[0] ? in[10] : in[9];
	assign out1[8] = shift[0] ? in[9] : in[8];
	assign out1[7] = shift[0] ? in[8] : in[7];
	assign out1[6] = shift[0] ? in[7] : in[6];
	assign out1[5] = shift[0] ? in[6] : in[5];
	assign out1[4] = shift[0] ? in[5] : in[4];
	assign out1[3] = shift[0] ? in[4] : in[3];
	assign out1[2] = shift[0] ? in[3] : in[2];
	assign out1[1] = shift[0] ? in[2] : in[1];
	assign out1[0] = shift[0] ? in[1] : in[0];
	
	// second layer 2
	assign out2[31] = shift[1] ? most_significant : out1[31];
	assign out2[30] = shift[1] ? most_significant : out1[30];
	assign out2[29] = shift[1] ? out1[31] : out1[29];
	assign out2[28] = shift[1] ? out1[30] : out1[28];
	assign out2[27] = shift[1] ? out1[29] : out1[27];
	assign out2[26] = shift[1] ? out1[28] : out1[26];
	assign out2[25] = shift[1] ? out1[27] : out1[25];
	assign out2[24] = shift[1] ? out1[26] : out1[24];
	assign out2[23] = shift[1] ? out1[25] : out1[23];
	assign out2[22] = shift[1] ? out1[24] : out1[22];
	assign out2[21] = shift[1] ? out1[23] : out1[21];
	assign out2[20] = shift[1] ? out1[22] : out1[20];
	assign out2[19] = shift[1] ? out1[21] : out1[19];
	assign out2[18] = shift[1] ? out1[20] : out1[18];
	assign out2[17] = shift[1] ? out1[19] : out1[17];
	assign out2[16] = shift[1] ? out1[18] : out1[16];
	assign out2[15] = shift[1] ? out1[17] : out1[15];
	assign out2[14] = shift[1] ? out1[16] : out1[14];
	assign out2[13] = shift[1] ? out1[15] : out1[13];
	assign out2[12] = shift[1] ? out1[14] : out1[12];
	assign out2[11] = shift[1] ? out1[13] : out1[11];
	assign out2[10] = shift[1] ? out1[12] : out1[10];
	assign out2[9] = shift[1] ? out1[11] : out1[9];
	assign out2[8] = shift[1] ? out1[10] : out1[8];
	assign out2[7] = shift[1] ? out1[9] : out1[7];
	assign out2[6] = shift[1] ? out1[8] : out1[6];
	assign out2[5] = shift[1] ? out1[7] : out1[5];
	assign out2[4] = shift[1] ? out1[6] : out1[4];
	assign out2[3] = shift[1] ? out1[5] : out1[3];
	assign out2[2] = shift[1] ? out1[4] : out1[2];
	assign out2[1] = shift[1] ? out1[3] : out1[1];
	assign out2[0] = shift[1] ? out1[2] : out1[0];
	
	
	// third layer 4
	assign out3[31] = shift[2] ? most_significant : out2[31];
	assign out3[30] = shift[2] ? most_significant : out2[30];
	assign out3[29] = shift[2] ? most_significant : out2[29];
	assign out3[28] = shift[2] ? most_significant : out2[28];
	assign out3[27] = shift[2] ? out2[31] : out2[27];
	assign out3[26] = shift[2] ? out2[30] : out2[26];
	assign out3[25] = shift[2] ? out2[29] : out2[25];
	assign out3[24] = shift[2] ? out2[28] : out2[24];
	assign out3[23] = shift[2] ? out2[27] : out2[23];
	assign out3[22] = shift[2] ? out2[26] : out2[22];
	assign out3[21] = shift[2] ? out2[25] : out2[21];
	assign out3[20] = shift[2] ? out2[24] : out2[20];
	assign out3[19] = shift[2] ? out2[23] : out2[19];
	assign out3[18] = shift[2] ? out2[22] : out2[18];
	assign out3[17] = shift[2] ? out2[21] : out2[17];
	assign out3[16] = shift[2] ? out2[20] : out2[16];
	assign out3[15] = shift[2] ? out2[19] : out2[15];
	assign out3[14] = shift[2] ? out2[18] : out2[14];
	assign out3[13] = shift[2] ? out2[17] : out2[13];
	assign out3[12] = shift[2] ? out2[16] : out2[12];
	assign out3[11] = shift[2] ? out2[15] : out2[11];
	assign out3[10] = shift[2] ? out2[14] : out2[10];
	assign out3[9] = shift[2] ? out2[13] : out2[9];
	assign out3[8] = shift[2] ? out2[12] : out2[8];
	assign out3[7] = shift[2] ? out2[11] : out2[7];
	assign out3[6] = shift[2] ? out2[10] : out2[6];
	assign out3[5] = shift[2] ? out2[9] : out2[5];
	assign out3[4] = shift[2] ? out2[8] : out2[4];
	assign out3[3] = shift[2] ? out2[7] : out2[3];
	assign out3[2] = shift[2] ? out2[6] : out2[2];
	assign out3[1] = shift[2] ? out2[5] : out2[1];
	assign out3[0] = shift[2] ? out2[4] : out2[0];
	
	// fourth layer 8
	assign out4[31] = shift[3] ? most_significant : out3[31];
	assign out4[30] = shift[3] ? most_significant : out3[30];
	assign out4[29] = shift[3] ? most_significant : out3[29];
	assign out4[28] = shift[3] ? most_significant : out3[28];
	assign out4[27] = shift[3] ? most_significant : out3[27];
	assign out4[26] = shift[3] ? most_significant : out3[26];
	assign out4[25] = shift[3] ? most_significant : out3[25];
	assign out4[24] = shift[3] ? most_significant : out3[24];
	assign out4[23] = shift[3] ? out3[31] : out3[23];
	assign out4[22] = shift[3] ? out3[30] : out3[22];
	assign out4[21] = shift[3] ? out3[29] : out3[21];
	assign out4[20] = shift[3] ? out3[28] : out3[20];
	assign out4[19] = shift[3] ? out3[27] : out3[19];
	assign out4[18] = shift[3] ? out3[26] : out3[18];
	assign out4[17] = shift[3] ? out3[25] : out3[17];
	assign out4[16] = shift[3] ? out3[24] : out3[16];
	assign out4[15] = shift[3] ? out3[23] : out3[15];
	assign out4[14] = shift[3] ? out3[22] : out3[14];
	assign out4[13] = shift[3] ? out3[21] : out3[13];
	assign out4[12] = shift[3] ? out3[20] : out3[12];
	assign out4[11] = shift[3] ? out3[19] : out3[11];
	assign out4[10] = shift[3] ? out3[18] : out3[10];
	assign out4[9] = shift[3] ? out3[17] : out3[9];
	assign out4[8] = shift[3] ? out3[16] : out3[8];
	assign out4[7] = shift[3] ? out3[15] : out3[7];
	assign out4[6] = shift[3] ? out3[14] : out3[6];
	assign out4[5] = shift[3] ? out3[13] : out3[5];
	assign out4[4] = shift[3] ? out3[12] : out3[4];
	assign out4[3] = shift[3] ? out3[11] : out3[3];
	assign out4[2] = shift[3] ? out3[10] : out3[2];
	assign out4[1] = shift[3] ? out3[9] : out3[1];
	assign out4[0] = shift[3] ? out3[8] : out3[0];
	
	
	// fifth layer 16
	assign out[31] = shift[4] ? most_significant : out4[31];
	assign out[30] = shift[4] ? most_significant : out4[30];
	assign out[29] = shift[4] ? most_significant : out4[29];
	assign out[28] = shift[4] ? most_significant : out4[28];
	assign out[27] = shift[4] ? most_significant : out4[27];
	assign out[26] = shift[4] ? most_significant : out4[26];
	assign out[25] = shift[4] ? most_significant : out4[25];
	assign out[24] = shift[4] ? most_significant : out4[24];
	assign out[23] = shift[4] ? most_significant : out4[23];
	assign out[22] = shift[4] ? most_significant : out4[22];
	assign out[21] = shift[4] ? most_significant : out4[21];
	assign out[20] = shift[4] ? most_significant : out4[20];
	assign out[19] = shift[4] ? most_significant : out4[19];
	assign out[18] = shift[4] ? most_significant : out4[18];
	assign out[17] = shift[4] ? most_significant : out4[17];
	assign out[16] = shift[4] ? most_significant : out4[16];
	assign out[15] = shift[4] ? out4[31] : out4[15];
	assign out[14] = shift[4] ? out4[30] : out4[14];
	assign out[13] = shift[4] ? out4[29] : out4[13];
	assign out[12] = shift[4] ? out4[28] : out4[12];
	assign out[11] = shift[4] ? out4[27] : out4[11];
	assign out[10] = shift[4] ? out4[26] : out4[10];
	assign out[9] = shift[4] ? out4[25] : out4[9];
	assign out[8] = shift[4] ? out4[24] : out4[8];
	assign out[7] = shift[4] ? out4[23] : out4[7];
	assign out[6] = shift[4] ? out4[22] : out4[6];
	assign out[5] = shift[4] ? out4[21] : out4[5];
	assign out[4] = shift[4] ? out4[20] : out4[4];
	assign out[3] = shift[4] ? out4[19] : out4[3];
	assign out[2] = shift[4] ? out4[18] : out4[2];
	assign out[1] = shift[4] ? out4[17] : out4[1];
	assign out[0] = shift[4] ? out4[16] : out4[0];
	
endmodule 